// -----------------------------------------------------------------------------
// Module: xorshift32 (Xorshift Pseudo-Random Number Generator)
// Author: MrAbhi19
// Description:
//   This module implements the Xorshift32 algorithm, a fast and lightweight
//   pseudo-random number generator based on XOR and bit-shift operations.
//
//   The generator evolves its internal 32-bit state on each clock cycle
//   (when enabled), producing a new pseudo-random number.
//
// Algorithm:
//   The recurrence relation is defined as:
//       X ^= (X << 13);
//       X ^= (X >> 17);
//       X ^= (X << 5);
//   where X is the internal state.
//
// Parameters:
//   None (constants are fixed for Xorshift32)
//
// Ports:
//   clk   - Input clock signal. Advances the generator on each rising edge.
//   rst   - Asynchronous reset. Resets the generator state to the seed.
//   en    - Enable signal. When high, the generator updates its state.
//   seed  - 32-bit input seed value used to initialize the generator.
//           Valid range: 1 to (2^32 - 1).
//   out   - 32-bit output representing the current pseudo-random number.
//
// Notes:
//   - Xorshift generators are known for speed and simplicity, but not for
//     cryptographic security. They are suitable for simulations, games,
//     and non-secure randomization tasks.
//   - The output sequence is deterministic given the same seed.
//   - Ensure the seed is non-zero to avoid a stuck state (all zeros).
// -----------------------------------------------------------------------------

module xorshift32 (
  input        clk,        // Clock input
  input        rst,        // Asynchronous reset input
  input        en,         // Enable input
  input  [31:0] seed,      // Seed value (1 to 2^32 - 1)
  output reg [31:0] out    // Current pseudo-random output
);

  reg [31:0] state;        // Internal state register

  // Sequential logic: update state and output on clock or reset
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      state <= seed;        // Initialize state with seed
      out   <= 0;           // Clear output on reset
    end else if (en) begin
      // Xorshift32 algorithm steps:
      state <= state ^ (state << 13); // Step 1: XOR with left shift by 13
      state <= state ^ (state >> 17); // Step 2: XOR with right shift by 17
      state <= state ^ (state << 5);  // Step 3: XOR with left shift by 5

      out   <= state;       // Update output with new state
    end
  end

endmodule
