// -----------------------------------------------------------------------------
// Module: lcg (Linear Congruential Generator)
// Author: MrAbhi19
// Description:
//   This module implements a simple Linear Congruential Generator (LCG),
//   which is a pseudo-random number generator defined by the recurrence:
//       X_{n+1} = (A * X_n + C) mod M
//
//   Each clock cycle produces the next pseudo-random number in the sequence.
//   The generator is initialized with a seed value.
//
// Parameters:
//   A - Multiplier constant (default = 214013)
//   C - Increment constant (default = 2531011)
//   M - Modulus constant (default = 2^31)
//
//  Microsoft C Runtime (MSVCRT) Variant:
//     - A = 214013
//     - C = 2531011
//     - M = 2^31
//     This is the widely used LCG configuration in Microsoft's C standard library.
//     Using these values will replicate the pseudo-random sequence generated by
//     the MSVCRT `rand()` function.
//
// Ports:
//   clk   - Input clock signal. Advances the generator on each rising edge.
//   rst   - Asynchronous reset. Resets the generator state to the seed.
//   seed  - 8-bit input seed value used to initialize the generator.
//   out   - 8-bit output representing the current pseudo-random number.
//
// Notes:
//   - The modulo operator (%) may not synthesize efficiently for non-power-of-2 M.
//     For hardware optimization, consider restricting M to powers of 2.
//   - This design is sequential and requires a clock for proper operation.
//   - The output sequence is deterministic given the same seed and parameters.
// -----------------------------------------------------------------------------

module lcg #(
  parameter A = 214013,   // Multiplier constant
  parameter C = 2531011,    // Increment constant
  parameter M = 2^31    // Modulus constant
)(
  input        clk,   // Clock input
  input        rst,   // Asynchronous reset input
  input  [7:0] seed,  // Seed value to initialize the generator
  output reg [7:0] out // Current pseudo-random output
);

  reg [7:0] inter;    // Internal state register

  // Sequential logic: update state and output on clock or reset
  always @(posedge clk or posedge rst) begin
    if (rst) begin
      inter <= seed;        // Initialize state with seed
      out   <= seed % M;    // Ensure output is within modulus range
    end else begin
      inter <= (inter * A + C) % M; // Compute next state
      out   <= inter;               // Update output
    end
  end

endmodule
